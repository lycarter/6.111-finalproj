`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:10:20 11/17/2016 
// Design Name: 
// Module Name:    debounce 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: Pushbutton Debounce Module (video version - 24 bits)  
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module debounce (input reset, clock, noisy,
                 output reg clean);

	reg [19:0] count;
    reg new;

    always @(posedge clock)
		if (reset) begin new <= noisy; clean <= noisy; count <= 0; end
		else if (noisy != new) begin new <= noisy; count <= 0; end
		else if (count == 650000) clean <= new;
		else count <= count+1;

endmodule
